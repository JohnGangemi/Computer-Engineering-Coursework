Inverter SPICE DECK				
**-----------------------------------------------------------------------------------------------------------------------
*   	Filename:	inverter.sp	
*	Author:		John Gangemi
*	Email:		JohnGangemi@mail.usf.edu
**-----------------------------------------------------------------------------------------------------------------------
* Parameters and models
**-----------------------------------------------------------------------------------------------------------------------
	.param SUPPLY = 5.0V            
   	.param GROUND = 0.0V		 
	.option post = ASCII 						
	.option list							 
	.option scale = 1u 						
	.option RUNLVL = 6			
	.temp 27							
	.lib '$USFCDK_HSPICE_PATH/SCN3ME_SUBM.lib' TT

**-----------------------------------------------------------------------------------------------------------------------
* Simulation Stimuli		
**-----------------------------------------------------------------------------------------------------------------------

 	Vdd    vdd    	gnd    'SUPPLY'

	.vec 'inverter.dat'

**-----------------------------------------------------------------------------------------------------------------------
* Simulation Netlist
**-----------------------------------------------------------------------------------------------------------------------

	.include netlist

**-----------------------------------------------------------------------------------------------------------------------
* Capacitive Loads
**-----------------------------------------------------------------------------------------------------------------------

	cl0 	z	gnd	0.01pF	

**-----------------------------------------------------------------------------------------------------------------------
* Parameters and models
**-----------------------------------------------------------------------------------------------------------------------
   
	.tran 0.1ns 30ns
	.print  tran V(a) V(z)

    .end
