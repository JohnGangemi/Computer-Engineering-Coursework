ThreeInputNOR SPICE DECK				* The first line is the title line of the simulation (max length is 72)
**-----------------------------------------------------------------------------------------------------------------------
*   	Filename:	ThreeInputNOR.sp	
*	Author: 	John A. Gangemi
*	Email:		JohnGangemi@mail.usf.edu
*	Class:		CDA4213L.F[14]
**-----------------------------------------------------------------------------------------------------------------------
* Parameters and models
**-----------------------------------------------------------------------------------------------------------------------
	.param SUPPLY = 5.0V            * 'SUPPLY' variable with value of 5.0V
   	.param GROUND = 0.0V		* 'GROUND' variable with value of 0.0V
	.param LOW = '(0.10*SUPPLY)'      * 'LOW' variable with value of 10% SUPPLY
	.param MID = '(0.50*SUPPLY)'     * 'MID' variable with value of 50% SUPPLY
	.param HIGH = '(0.90*SUPPLY)'     * 'HIGH' variable with value of 90% SUPPLY
	.option post = ASCII 						
	.option list							 
	.option scale = 1u 						
	.option RUNLVL = 6			
	.temp 27	
	.lib '$USFCDK_HSPICE_PATH/SCN3ME_SUBM.lib' TT							

**-----------------------------------------------------------------------------------------------------------------------
* Simulation Stimuli
**-----------------------------------------------------------------------------------------------------------------------
*
*	V[id]  N1	  gnd	 Value	
*
**-----------------------------------------------------------------------------------------------------------------------
    Vdd    vdd    gnd    'SUPPLY'

    **********************************************************
    ** Uncomment labeled sections to test different stimuli **
    ** Vector data is default and therefore uncommented     **
    **********************************************************

    * PULSE INPUT STIMULI *
    ***********************

    *VA    A      gnd	 PULSE 'GROUND' 'SUPPLY' 0.0ns 0.1ns 0.1ns 15ns 30ns
    *VB	   B	  gnd	 PULSE 'GROUND' 'SUPPLY' 0.0ns 0.1ns 0.1ns 5ns 10ns
    *VC	   C	  gnd	 PULSE 'GROUND' 'SUPPLY' 0.0ns 0.1ns 0.1ns 5ns 10ns

    * VECTOR INPUT STIMULI *
    ************************

    .vec 'ThreeInputNOR.dat'
		
**-----------------------------------------------------------------------------------------------------------------------
*
*	PULSE 'Low Voltage' 'High Voltage' 'StartTime' 'RiseTime' 'FallTime' 'TimeHigh' 'TotalCycle'
*
*	PWL 'TimeX' 'VoltageX' 'TimeX+1' 'VoltageX+1' ....... 'TimeN' 'VoltageN'
*
**-----------------------------------------------------------------------------------------------------------------------
* Simulation Netlist
**-----------------------------------------------------------------------------------------------------------------------
	.include ThreeInputNORnetlist		* Includes the content of the specified file 'netlist'
**-----------------------------------------------------------------------------------------------------------------------	
*
*	C[id]  N1     N2    Value	 <IC>		* Generic format for cload statements
*
**-----------------------------------------------------------------------------------------------------------------------
	cl0    Z     gnd   0.01pF
**-----------------------------------------------------------------------------------------------------------------------
* Stimulus
**-----------------------------------------------------------------------------------------------------------------------
*
*	.tran	Interval	StopTime
*
**-----------------------------------------------------------------------------------------------------------------------
	.tran   0.1ns 80ns			 * Performs and prints the transient analysis, every .1 ns for 80 ns

**-----------------------------------------------------------------------------------------------------------------------
* Parameters and models
**-----------------------------------------------------------------------------------------------------------------------
*
*	.print	tran   V(in0) V(in1) ...... V(out0) V(out1)......
*
**-----------------------------------------------------------------------------------------------------------------------    
	.print  tran V(A) V(B) V(C) V(Z)

**-----------------------------------------------------------------------------------------------------------------------
* Alterations / Resimulations
**-----------------------------------------------------------------------------------------------------------------------
	
**-----------------------------------------------------------------------------------------------------------------------
* EOF
**-----------------------------------------------------------------------------------------------------------------------
    .end
